library IEEE;use IEEE.STD_LOGIC_1164.ALL;use IEEE.STD_LOGIC_ARITH.ALL;use IEEE.STD_LOGIC_UNSIGNED.ALL;library work;--use work.adcmv3_components.all;entity shower_spi_adc_master isgeneric(	RESET_VALUE_CTRL    : std_logic_vector(7 downto 0) := x"00");port(CLK_IN          : in    std_logic;	RESET_IN        : in    std_logic;	-- Slave bus	SLV_READ_IN     : in    std_logic;	SLV_WRITE_IN    : in    std_logic;	SLV_BUSY_OUT    : out   std_logic;	SLV_ACK_OUT     : out   std_logic;	SLV_DATA_IN     : in    std_logic_vector(31 downto 0);	SLV_DATA_OUT    : out   std_logic_vector(31 downto 0);	-- SPI connections	SPI_CS_OUT      : out   std_logic;	SPI_SDO_OUT     : out   std_logic;	SPI_SCK_OUT     : out   std_logic;	-- ADC connections	ADC_LOCKED_IN   : in    std_logic;	ADC_PD_OUT      : out   std_logic;	ADC_RST_OUT     : out   std_logic;	ADC_DEL_OUT     : out   std_logic_vector(3 downto 0);	-- Status lines	STAT            : out   std_logic_vector(31 downto 0) -- DEBUG);end entity;architecture Behavioral of shower_spi_adc_master is-- Componentscomponent shower_spi_real_slim isport(	SYSCLK      : in    std_logic; -- 100MHz sysclock	RESET       : in    std_logic; -- synchronous reset	-- Command interface	START_IN    : in    std_logic; -- one start pulse	BUSY_OUT    : out   std_logic; -- SPI transactions are ongoing	CMD_IN      : in    std_logic_vector(23 downto 0); -- SPI command byte	-- SPI interface	SPI_SCK_OUT : out   std_logic;	SPI_CS_OUT  : out   std_logic;	SPI_SDO_OUT : out   std_logic;	-- DEBUG	CLK_EN_OUT  : out   std_logic;	BSM_OUT     : out   std_logic_vector(7 downto 0);	DEBUG_OUT   : out   std_logic_vector(31 downto 0));end component shower_spi_real_slim;-- Signalstype STATES is (SLEEP,RD_BSY,WR_BSY,RD_RDY,WR_RDY,RD_ACK,WR_ACK,DONE);signal CURRENT_STATE, NEXT_STATE: STATES;signal status_data      : std_logic_vector(31 downto 0);signal spi_busy         : std_logic;signal reg_ctrl_data    : std_logic_vector(23 downto 0);signal adc_ctrl_data    : std_logic_vector(7 downto 0);signal reg_slv_data_out : std_logic_vector(31 downto 0); -- readbacksignal spi_start_x      : std_logic;signal spi_start        : std_logic;-- State machine signalssignal slv_busy_x       : std_logic;signal slv_busy         : std_logic;signal slv_ack_x        : std_logic;signal slv_ack          : std_logic;signal store_wr_x       : std_logic;signal store_wr         : std_logic;signal store_rd_x       : std_logic;signal store_rd         : std_logic;begin----------------------------------------------------------- SPI master                                          -----------------------------------------------------------THE_SPI_REAL_SLIM: shower_spi_real_slimport map(	SYSCLK      => clk_in,	RESET       => reset_in,	-- Command interface	START_IN    => spi_start,	BUSY_OUT    => spi_busy,	CMD_IN      => reg_ctrl_data,	-- SPI interface	SPI_SCK_OUT => spi_sck_out,	SPI_CS_OUT  => spi_cs_out,	SPI_SDO_OUT => spi_sdo_out,	-- DEBUG	CLK_EN_OUT  => open,	BSM_OUT     => open,	DEBUG_OUT   => open);----------------------------------------------------------- Statemachine                                        ------------------------------------------------------------- State memory processSTATE_MEM: process( clk_in )begin	if( rising_edge(clk_in) ) then		if( reset_in = '1' ) then			CURRENT_STATE <= SLEEP;			slv_busy      <= '0';			slv_ack       <= '0';			store_wr      <= '0';			store_rd      <= '0';		else			CURRENT_STATE <= NEXT_STATE;			slv_busy      <= slv_busy_x;			slv_ack       <= slv_ack_x;			store_wr      <= store_wr_x;			store_rd      <= store_rd_x;		end if;	end if;end process STATE_MEM;-- Transition matrixTRANSFORM: process(CURRENT_STATE, slv_read_in, slv_write_in, spi_busy )begin	NEXT_STATE <= SLEEP;	slv_busy_x <= '0';	slv_ack_x  <= '0';	store_wr_x <= '0';	store_rd_x <= '0';	case CURRENT_STATE is		when SLEEP      =>  if   ( (spi_busy = '0') and (slv_read_in = '1') ) then								NEXT_STATE <= RD_RDY;								store_rd_x <= '1';							elsif( (spi_busy = '0') and (slv_write_in = '1') ) then								NEXT_STATE <= WR_RDY;								store_wr_x <= '1';							elsif( (spi_busy = '1') and (slv_read_in = '1') ) then								NEXT_STATE <= RD_BSY;								slv_busy_x <= '1';							elsif( (spi_busy = '1') and (slv_write_in = '1') ) then								NEXT_STATE <= WR_BSY;								slv_busy_x <= '1';							else								NEXT_STATE <= SLEEP;							end if;		when RD_RDY     =>  NEXT_STATE <= RD_ACK;							slv_ack_x  <= '1';		when WR_RDY     =>  NEXT_STATE <= WR_ACK;							slv_ack_x  <= '1';		when RD_ACK     =>  if( slv_read_in = '0' ) then								NEXT_STATE <= DONE;							else								NEXT_STATE <= RD_ACK;								slv_ack_x  <= '1';							end if;		when WR_ACK     =>  if( slv_write_in = '0' ) then								NEXT_STATE <= DONE;							else								NEXT_STATE <= WR_ACK;								slv_ack_x  <= '1';							end if;		when RD_BSY     =>  if( slv_read_in = '0' ) then								NEXT_STATE <= DONE;							else								NEXT_STATE <= RD_BSY;								slv_busy_x <= '1';							end if;		when WR_BSY     =>  if( slv_write_in = '0' ) then								NEXT_STATE <= DONE;							else								NEXT_STATE <= WR_BSY;								slv_busy_x <= '1';							end if;		when DONE       =>  NEXT_STATE <= SLEEP;		when others     =>  NEXT_STATE <= SLEEP;	end case;end process TRANSFORM;----------------------------------------------------------- data handling                                       ------------------------------------------------------------- register writeTHE_WRITE_REG_PROC: process( clk_in )begin	if( rising_edge(clk_in) ) then		if   ( reset_in = '1' ) then			reg_ctrl_data   <= (others => '0');			adc_ctrl_data   <= RESET_VALUE_CTRL;			spi_start       <= '0';		elsif( store_wr = '1' ) then			reg_ctrl_data   <= slv_data_in(31 downto 8 );			adc_ctrl_data   <= slv_data_in(7 downto 0);		end if;		spi_start <= spi_start_x;	end if;end process THE_WRITE_REG_PROC;spi_start_x <= '1' when ( (store_wr = '1') and (slv_data_in(3) = '1') ) else '0';-- register readTHE_READ_REG_PROC: process( clk_in )begin	if( rising_edge(clk_in) ) then		if   ( reset_in = '1' ) then			reg_slv_data_out <= (others => '0');		elsif( store_rd = '1' ) then			reg_slv_data_out <= reg_ctrl_data & adc_ctrl_data;		end if;	end if;end process THE_READ_REG_PROC;-- debug signalsstatus_data(31 downto 0)  <= (others => '0');-- output signalsadc_del_out  <= adc_ctrl_data(7 downto 4);adc_pd_out   <= adc_ctrl_data(1);adc_rst_out  <= not adc_ctrl_data(0);stat         <= status_data;slv_ack_out  <= slv_ack;slv_busy_out <= slv_busy;slv_data_out <= reg_slv_data_out;end Behavioral;
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:19:23 09/27/2008 
-- Design Name: 
-- Module Name:    read_ADCs - Behavioral 
-- Project Name: 

-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- use IEEE.STD_LOGIC_ARITH.ALL;
-- use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.numeric_std.all;
use work.shower_components.all;

entity read_ADC is
       generic (
         IOFF_DELAY   : std_logic_vector(3 downto 0) :=  "0000"
         );

    port (  RESET         : in std_logic;
      CLOCK         : in std_logic; 
--         --Pedestal / connection to bus handler
    PED_DATA_IN            : in std_logic_vector(9 downto 0);
    PED_DATA_OUT           : out std_logic_vector(9 downto 0);
        TRB_PED_ADDR_IN        : in std_logic_vector(8 downto 0);
        PED_READ_IN            : in std_logic;
        PED_WRITE_IN           : in std_logic;
        PED_READ_ACK_OUT       : out std_logic;
        PED_WRITE_ACK_OUT      : out std_logic;
        PED_BUSY_OUT           : out std_logic;
        PED_UNKNOWN_OUT        : out std_logic;
  
      IOFF_DELAY_IN     : in std_logic_vector(3 downto 0);
      LOCAL_ID_IN       : in std_logic_vector(3 downto 0);
      SAMPLING_PATTERN_IN   : in std_logic_vector (3 downto 0);
      THRESHOLD_IN      : in std_logic_vector (3 downto 0);

         --ADC inputs
      ADC_DATA_CLOCK_IN       : in std_logic;
      ADC_FRAME_CLOCK_IN      : in std_logic;
      ADC_SERIAL_IN   : in std_logic_vector(7 downto 0);

--         --Control signals from FEB
-- 10 ns pulse when FEB multiplexer advances input channel
      FEB_MUX_NEW_CHAN_RDY_IN : in std_logic;
      FEB_64TH_PEDESTAL_OUT : out std_logic;
      --  data interface to endpint handler
      FEE_TRG_TYPE_IN     : in std_logic_vector(3  downto 0);
      FEE_TRG_DATA_VALID_IN  :   in std_logic;
      FEE_DATA_OUT      : out std_logic_vector(31 downto 0);
      FEE_DATA_WRITE_OUT    : out std_logic;
      FEE_DATA_FINISHED_OUT : out std_logic;

         --Data Output to ipu_han
        IPU_DAT_DATA_OUT      : out std_logic_vector(26 downto 0);
        IPU_DAT_DATA_READ_IN  : in std_logic;
        IPU_DAT_DATA_EMPTY_OUT : out std_logic;
        IPU_HDR_DATA_OUT      : out std_logic_vector(17 downto 0);
        IPU_HDR_DATA_READ_IN  : in std_logic;
        IPU_HDR_DATA_EMPTY_OUT : out std_logic;
-- outputs to trb Slow Control REGIO_STAT_REG
        SERPAR_INPUT_FIFO_EMPTY :out std_logic;
        SERPAR_INPUT_FIFO_FULL  :out std_logic;
       --Debug
      ADC_INSPECT_BUS     : out std_logic_vector(35 downto 0));
end read_ADC;

architecture Behavioral of read_ADC is
--attribute HGROUP : string;
--attribute HGROUP of Behavioral : architecture is "ADC_chip";

type ADC_INPUT_VECTOR_ARRAY is array (7 downto 0) of std_logic_vector(0 downto 0);
type ADC_CHANN_ARRAY_12BIT is array (8 downto 1) of unsigned (11 downto 0);

type write_state_type is (idle, wait_for_average, wait_for_comparators, wait_for_comp_status, write_to_fifo, 
              inc_channel_counter, test_completed, column_finished, test_event_finished,
              event_finished, send_out_thresholds, event_finished_or_continue_pedestal);
--********************** MK
type PEDESTAL_DATA_ARRAY is array (8 downto 1) of unsigned (15 downto 0);

type acalcul_state_type is (idle_ac, first_pedestal_sample, write_ADC_to_memory, check_first_event_end,
check_counter, wait_for_next_event, read_pedestal_value, sum_with_ADC, write_sum_to_memory,
check_ped_event_end, average_calcul_finished, synch_wait, synch_wait_1);

signal acalcul_state, next_acalcul_state : acalcul_state_type;
--********************** MK end

signal write_state, next_write_state : write_state_type;

attribute syn_encoding: string;
attribute syn_encoding of write_state: signal is "safe,onehot";

signal COLUMN_COUNTER : unsigned (10 downto 0);
signal PEDESTAL_ADDRESS : std_logic_vector(4 downto 0);
signal WIDE_ADC_BUS  : std_logic_vector(79 downto 0);
--signal WIDER_ADC_BUS  : unsigned(95 downto 0);
signal ADC_IN_BUS : std_logic_vector(9 downto 0);
signal ADC_THRESHOLD_BUS : std_logic_vector(9 downto 0);
signal channel_threshold : PEDESTAL_OUT_ARRAY;
signal WRITE_PEDESTAL : std_logic_vector(8 downto 1);
signal ADC_INPUT_VECTOR     : ADC_INPUT_VECTOR_ARRAY;
signal ADC_INPUT_7, ADC_INPUT_6, ADC_INPUT_5, ADC_INPUT_4 : std_logic_vector(0 downto 0);
signal ADC_INPUT_3, ADC_INPUT_2, ADC_INPUT_1, ADC_INPUT_0 : std_logic_vector(0 downto 0);
signal FRAME_CLOCK_VECTOR : std_logic_vector(0 downto 0);
signal sampled_FRAME_CLOCK : std_logic_vector(1 downto 0);
signal sampled_ADC_INPUT : std_logic_vector(15 downto 0);
signal execute_write : std_logic;
signal ADC_RESULT_VALID, serpar_full, serpar_empty : std_logic;

signal integrator, average : ADC_CHANN_ARRAY_12BIT; 

signal sampling_end : std_logic_vector (7 downto 0);
signal current_sampling_pattern : std_logic_vector (5 downto 0);
signal delayed_start : std_logic_vector (8 downto 0);
signal start_extended: std_logic;
signal channel_counter : unsigned (3 downto 0);
signal comp_result, threshold_comparison_status : std_logic_vector (7 downto 0);
signal add_result : std_logic_vector (95 downto 0);

signal inverted_sampling_pattern : std_logic_vector (0 to 3);
signal fee_trg_type: std_logic_vector(3  downto 0);
signal fee_data_finished : std_logic;
signal fee_data_write : std_logic;

signal pedestal_calculation : std_logic;
signal PEDESTAL_DATA_IN_16, pedestal_sum : PEDESTAL_DATA_ARRAY;
signal PEDESTAL_EVENT_COUNTER : unsigned (5 downto 0);

signal state_bits: std_logic_vector(3 downto 0);
signal SERPAR_INSPECT_BUS: std_logic_vector(31 downto 0);

signal delayed_write_ack, delayed_read_ack : std_logic_vector(2 downto 0);

attribute syn_preserve : boolean;
attribute syn_preserve of write_state : signal is true;
attribute syn_preserve of COLUMN_COUNTER : signal is true;

begin

FEE_DATA_FINISHED_OUT <= fee_data_finished;
FEE_DATA_WRITE_OUT <= fee_data_write;
FRAME_CLOCK_VECTOR(0) <= ADC_FRAME_CLOCK_IN;

ADC_INPUT_7(0) <= ADC_SERIAL_IN(7);
ADC_INPUT_6(0) <= ADC_SERIAL_IN(6);
ADC_INPUT_5(0) <= ADC_SERIAL_IN(5);
ADC_INPUT_4(0) <= ADC_SERIAL_IN(4);
ADC_INPUT_3(0) <= ADC_SERIAL_IN(3);
ADC_INPUT_2(0) <= ADC_SERIAL_IN(2);
ADC_INPUT_1(0) <= ADC_SERIAL_IN(1);
ADC_INPUT_0(0) <= ADC_SERIAL_IN(0);

-- modelssim display file : draw_adc-simple1
--ADC_INSPECT_BUS <= '0' &  
--            sampling_end(4) & 
--            current_sampling_pattern(5) &
--            threshold_comparison_status(1 downto 0) & 
--            channel_counter(2 downto 0) & 
--            average(9 downto 0) &
--            FEE_DATA_WRITE_OUT & 
--            ADC_RESULT_VALID & 
--            delayed_start(8) & 
--            FEE_DATA_FINISHED_OUT &
--            channel_threshold(1);

ADC_INSPECT_BUS <= x"0000000" & delayed_start(8) & sampling_end(5) & start_extended & ADC_RESULT_VALID & SERPAR_INSPECT_BUS(23 downto 20);
--ADC_INSPECT_BUS <= SERPAR_INSPECT_BUS(31 downto 4) & state_bits;
--ADC_INSPECT_BUS <= sampled_FRAME_CLOCK & sampled_ADC_INPUT & SERPAR_INSPECT_BUS(17 downto 0);

-- THE_ADC_HANDLER : shower_adc_data_handler
--         port map(
--             CLK_IN => CLOCK,                    -- SYSCLK from fabric
--             RESET_IN => RESET,                  -- synchronous reset (SYSCLK clock domain)
--             ADC_RESET_IN => '0',
-- 
--             ADC_DCO_IN => ADC_DATA_CLOCK_IN,   -- DCO clock from ADC (direct I/O connection)
--             ADC_FCO_IN => ADC_FRAME_CLOCK_IN, -- FCO clock from ADC (direct I/O connection)
--             ADC_CHNL_IN => ADC_SERIAL_IN,       -- DDR data stream from ADC (direct I/O connection)
-- 
--             ADC_DATA7_OUT => WIDE_ADC_BUS(79 downto 70), -- parallel ADC data stream (7)
--             ADC_DATA6_OUT => WIDE_ADC_BUS(69 downto 60), -- parallel ADC data stream (6)
--             ADC_DATA5_OUT => WIDE_ADC_BUS(59 downto 50), -- parallel ADC data stream (5)
--             ADC_DATA4_OUT => WIDE_ADC_BUS(49 downto 40), -- parallel ADC data stream (4)
--             ADC_DATA3_OUT => WIDE_ADC_BUS(39 downto 30), -- parallel ADC data stream (3)
--             ADC_DATA2_OUT => WIDE_ADC_BUS(29 downto 20), -- parallel ADC data stream (2)
--             ADC_DATA1_OUT => WIDE_ADC_BUS(19 downto 10), -- parallel ADC data stream (1)
--             ADC_DATA0_OUT => WIDE_ADC_BUS( 9 downto  0), -- parallel ADC data stream (0)
-- 
--             ADC_CE_OUT => ADC_RESULT_VALID,              -- ADC data valid signal, centered into valid data
-- 
--             DEBUG_OUT =>  SERPAR_INSPECT_BUS(15 downto 0)
--         );

  THE_FCLK_DDR_FF : ddr_input_ff --ddr_iff_sysclk 
        port map(
            Del  => "0000",
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => FRAME_CLOCK_VECTOR,
            Q    => sampled_FRAME_CLOCK
            );

  THE_DATA_DDR_FF_0 : ddr_input_ff --ddr_iff_sysclk  
        port map(
            Del  => IOFF_DELAY_IN,
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => ADC_INPUT_0,
            Q(0)    => sampled_ADC_INPUT(1),
            Q(1)    => sampled_ADC_INPUT(0)
            );
  THE_DATA_DDR_FF_1 : ddr_input_ff --ddr_iff_sysclk  
        port map(
            Del  => IOFF_DELAY_IN,  
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => ADC_INPUT_1,
            Q(0)    => sampled_ADC_INPUT(3),
            Q(1)    => sampled_ADC_INPUT(2)
            );
  THE_DATA_DDR_FF_2 : ddr_input_ff --ddr_iff_sysclk  
        port map(
            Del  => IOFF_DELAY_IN,
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => ADC_INPUT_2,
            Q(0)    => sampled_ADC_INPUT(5),
            Q(1)    => sampled_ADC_INPUT(4)
            );
  THE_DATA_DDR_FF_3 : ddr_input_ff --ddr_iff_sysclk  
        port map(
            Del  => IOFF_DELAY_IN,
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => ADC_INPUT_3,
            Q(0)    => sampled_ADC_INPUT(7),
            Q(1)    => sampled_ADC_INPUT(6)
            );
  THE_DATA_DDR_FF_4 : ddr_input_ff --ddr_iff_sysclk  
        port map(
            Del  => IOFF_DELAY_IN,
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => ADC_INPUT_4,
            Q(0)    => sampled_ADC_INPUT(9),
            Q(1)    => sampled_ADC_INPUT(8)
            );
  THE_DATA_DDR_FF_5 : ddr_input_ff --ddr_iff_sysclk  
        port map(
            Del  => IOFF_DELAY_IN,
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => ADC_INPUT_5,
            Q(0)    => sampled_ADC_INPUT(11),
            Q(1)    => sampled_ADC_INPUT(10)
            );
  THE_DATA_DDR_FF_6 : ddr_input_ff --ddr_iff_sysclk  
        port map(
            Del  => IOFF_DELAY_IN,
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => ADC_INPUT_6,
            Q(0)    => sampled_ADC_INPUT(13),
            Q(1)    => sampled_ADC_INPUT(12)
            );
  THE_DATA_DDR_FF_7 : ddr_input_ff --ddr_iff_sysclk  
        port map(
            Del  => IOFF_DELAY_IN,
            CLK  => ADC_DATA_CLOCK_IN, --ECLK  => ADC_DATA_CLOCK_IN,
            --SCLK => CLOCK,
            Rst  => RESET,
            Data => ADC_INPUT_7,
            Q(0)    => sampled_ADC_INPUT(15),
            Q(1)    => sampled_ADC_INPUT(14)
            );

ADC: serpar2 port map (
    RESET         => RESET,
    ADC_CLOCK       => ADC_DATA_CLOCK_IN,
    SYS_CLOCK       => CLOCK,
    ADC_INPUT       => sampled_ADC_INPUT,
    FRAME_CLOCK     => sampled_FRAME_CLOCK,
    ADC_RESULT_OUT    => WIDE_ADC_BUS,
    ADC_RESULT_VALID_OUT  => ADC_RESULT_VALID,
      fifo_full       => SERPAR_INPUT_FIFO_FULL,
      fifo_empty      => SERPAR_INPUT_FIFO_EMPTY,
    debug             => SERPAR_INSPECT_BUS
    );

pedestal_memory: for i in 1 to 8 generate
pedestals: pedestal_DPRAM_32x16 port map (
  WrAddress   => PEDESTAL_ADDRESS,
  RdAddress   => PEDESTAL_ADDRESS,
  DATA      => std_logic_vector(PEDESTAL_DATA_IN_16(i)),
  WE        => WRITE_PEDESTAL(i),
  RdClock     => CLOCK,
  RdClockEn   => '1',
  Reset     => RESET,
    WrClock     => CLOCK,
  WrClockEn   => '1',
  Q       => channel_threshold(i));
end generate;

FEE_DATA_FINISHED_PROCESS: process (RESET, CLOCK, write_state) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    fee_data_finished <= '0';
  else
    if write_state = event_finished then
      fee_data_finished <= '1';
    else
      fee_data_finished <= '0';
    end if;
  end if;
end if; 
end process FEE_DATA_FINISHED_PROCESS;

FEE_TRG_TYPE_VALID_PROCESS: process (RESET, CLOCK, FEE_TRG_DATA_VALID_IN) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    fee_trg_type <= (others => '0');
  else
    if FEE_TRG_DATA_VALID_IN = '1' then
      fee_trg_type <= FEE_TRG_TYPE_IN;
    end if;
  end if;
end if; 
end process FEE_TRG_TYPE_VALID_PROCESS;

  
THR_COMPARISON_PROCESS: process(CLOCK, fee_trg_type) begin
if rising_edge(CLOCK) then
    if (fee_trg_type = x"A") or (fee_trg_type = x"B") then
    threshold_comparison_status <= "11111111";
  else 
    if write_state = wait_for_comp_status then 
      gen_test: for i in 0 to 7 loop
        if average(i+1)(9 downto 0) > (unsigned (channel_threshold(i+1)(15 downto 6)) + unsigned (THRESHOLD_IN)) then
          threshold_comparison_status(i) <= '1';
        else
          threshold_comparison_status(i) <= '0';
        end if;
      end loop;
    elsif write_state = test_completed then
        threshold_comparison_status <= '0' & threshold_comparison_status(7 downto 1);
    end if;
  end if;
end if;
end process THR_COMPARISON_PROCESS;

START_EXTENDED_PROCESS: process (RESET, CLOCK, FEB_MUX_NEW_CHAN_RDY_IN) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    start_extended <= '0';
  else
    if start_extended = '0' then
      if FEB_MUX_NEW_CHAN_RDY_IN = '1' then
        start_extended <= '1';
      end if;
    else
      if (delayed_start(0) = '1') then 
          start_extended <= '0';
      end if;
    end if;
  end if;
end if; 
end process START_EXTENDED_PROCESS;

--********************** MK

START_PEDEST_CAL_PROCESS: process (RESET, CLOCK, fee_trg_type) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    pedestal_calculation <= '0';
  else
    if pedestal_calculation = '0' then
      if fee_trg_type = x"B" and FEE_TRG_DATA_VALID_IN = '1' then
        pedestal_calculation <= '1';
      end if;
    else
      if write_state = event_finished then 
          pedestal_calculation <= '0';
      end if;
    end if;
  end if;
end if; 
end process START_PEDEST_CAL_PROCESS;

SELECT_PEDESTL_MEM_INPUT: process (RESET, CLOCK, acalcul_state) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    for i in 1 to 8 loop
      PEDESTAL_DATA_IN_16(i) <= unsigned(PED_DATA_IN & "000000");
    end loop;
  else
    if COLUMN_COUNTER(10 downto 5) = "000000" then
          gener_2 : for i in 1 to 8  loop
            PEDESTAL_DATA_IN_16(i) <= unsigned("0000" & average(i));
          end loop;
    else
          gener_3 : for i in 1 to 8  loop
            PEDESTAL_DATA_IN_16(i) <= pedestal_sum(i);
          end loop;
    end if;
 end if;
end if;
end process SELECT_PEDESTL_MEM_INPUT;

SUMMING_PEDESTAL: process (RESET, CLOCK) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    for i in 0 to 7 loop
      pedestal_sum(i+1) <= (others => '0');
    end loop;
  elsif write_state = wait_for_comparators then     --*******************
    gen_sum: for i in 0 to 7 loop
      pedestal_sum(i+1) <= unsigned(channel_threshold(i+1)) + unsigned("0000" & average(i+1));
    end loop;
  end if;
end if;
end process SUMMING_PEDESTAL;

COUNT_PED_TRIGGERS: process(RESET, CLOCK, write_state, acalcul_state) begin
if rising_edge(CLOCK) then
  if (RESET = '1') then
    PEDESTAL_EVENT_COUNTER <= (others => '0');
  else
    if write_state = event_finished and pedestal_calculation = '1' then   --******************
      PEDESTAL_EVENT_COUNTER <= PEDESTAL_EVENT_COUNTER + 1;
    else
      if acalcul_state = average_calcul_finished then
        PEDESTAL_EVENT_COUNTER <= (others => '0');
      end if;
    end if;
  end if;
end if;
end process COUNT_PED_TRIGGERS;

LAST_PEDESTAL: process (RESET, CLOCK, PEDESTAL_EVENT_COUNTER) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
      FEB_64TH_PEDESTAL_OUT <= '0';
  elsif PEDESTAL_EVENT_COUNTER = "111111" then
      FEB_64TH_PEDESTAL_OUT <= '1';
    else
      FEB_64TH_PEDESTAL_OUT <= '0';
  end if;
end if;
end process LAST_PEDESTAL;



SIMULATE_ADC_PIPE: process (RESET, CLOCK, ADC_RESULT_VALID) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    sampling_end <= (others => '0');
  else
    if (ADC_RESULT_VALID = '1') then             -- register shifts synchronously with ADC results (20 MSPS: every 50 ns)
      sampling_end <= sampling_end (6 downto 0) & delayed_start(7);  -- kk (8)
    end if;
  end if;
end if;
end process SIMULATE_ADC_PIPE;

DELAYED_COLUMN_PROCESS: process (RESET, CLOCK, ADC_RESULT_VALID) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    delayed_start <= (others => '0');
  else
    if (ADC_RESULT_VALID = '1') then             -- register shifts synchronously with ADC results (20 MSPS: every 50 ns)
      delayed_start <= delayed_start (7 downto 0) & start_extended;
    end if;
  end if;
end if;
end process DELAYED_COLUMN_PROCESS;

--inverted_sampling_pattern <= SAMPLING_PATTERN_IN;

MARK_VALID_SAMPLES_PROCESS: process (RESET, CLOCK) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    current_sampling_pattern <= "000000";
  else
    if ADC_RESULT_VALID = '1' then 
      if (delayed_start(6) = '1') then -- kk (8)
        current_sampling_pattern <= '0' &  SAMPLING_PATTERN_IN & '0';
      else
        current_sampling_pattern <= current_sampling_pattern (4 downto 0) & '0';
      end if;
    end if;
  end if;
end if;   
end process MARK_VALID_SAMPLES_PROCESS;

INTEGRATE_ADC_RESULTS_PROCESS: process (RESET, CLOCK) begin
if rising_edge (CLOCK) then
  if (RESET = '1' or write_state = wait_for_comparators) then -- reset integrator one clk after it has been copied to average
    for i in 1 to 8 loop
      integrator(i) <= (others => '0');
    end loop;
  else
    if ADC_RESULT_VALID = '1' and current_sampling_pattern(5) = '1' then
           gen_sum: for i in 0 to 7 loop
        integrator(i+1) <= integrator(i+1) + unsigned("00" & WIDE_ADC_BUS(10*i+9 downto 10*i));
            end loop;
        end if;
    end if;
end if;   
end process INTEGRATE_ADC_RESULTS_PROCESS;

AVERAGE_ADC_RESULTS_PROCESS: process (RESET, CLOCK) begin
if rising_edge (CLOCK) then
  if (RESET = '1') then
    for i in 1 to 8 loop
      average(i) <= (others => '0');
    end loop;
  else
    if write_state = wait_for_average then
        case SAMPLING_PATTERN_IN is
        when "0001"|"0010"|"0100"|"1000" =>     -- no division
          gen_div_1 : for i in 1 to 8 loop
            average(i) <= integrator (i);
          end loop;
        when "0011"|"0110"|"1100"|"1010"|"0101"|"1001" =>   -- division by 2 (shift by one bit)
          gen_div_2 : for i in 1 to 8 loop
            average(i) <= integrator (i) / 2;
          end loop;
        when "1111" =>                  -- division by 4 (shift by two bits)
          gen_div_4 : for i in 1 to 8 loop
            average(i) <= integrator (i) / 4;
          end loop;
        when others =>
          gen_div_1_others : for i in 1 to 8 loop
            average(i) <= integrator (i);
          end loop;
      end case;
        end if;
    end if;
end if;   
end process AVERAGE_ADC_RESULTS_PROCESS;

CHANNEL_COUNTER_PROCESS: process (RESET, CLOCK, write_state) begin
if rising_edge (CLOCK) then
  if (RESET = '1' or write_state = idle) then
    channel_counter <= (others =>'0');
  elsif write_state = write_to_fifo then
    channel_counter <= channel_counter + 1;
  end if;
end if;
end process CHANNEL_COUNTER_PROCESS;

ADC_IN_BUS_CC_PROC: process (RESET, CLOCK) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    FEE_DATA_OUT <= (others => '0');
  else
    if pedestal_calculation = '0' then
          FEE_DATA_OUT <= "000000000" & std_logic_vector(channel_counter (2 downto 0)) 
                        & "000" & std_logic_vector(COLUMN_COUNTER(4 downto 0)) & "00" & ADC_IN_BUS;
    else
          FEE_DATA_OUT <= "000000000" & std_logic_vector(channel_counter (2 downto 0)) 
                        & "000" & std_logic_vector(COLUMN_COUNTER(4 downto 0)) & "00" & ADC_IN_BUS;
    end if;
  end if;
end if;
end process ADC_IN_BUS_CC_PROC;

ADC_THRESHOLD_BUS_PROC: process (RESET, channel_counter)  begin
--if  rising_edge(CLOCK) then
  if (RESET = '1') then
  ADC_THRESHOLD_BUS <= (others => '0');
  else
  case std_logic_vector(channel_counter(2 downto 0)) is
    when "000"    => ADC_THRESHOLD_BUS <=  channel_threshold(1);
    when "001"    => ADC_THRESHOLD_BUS <=  channel_threshold(2);
    when "010"    => ADC_THRESHOLD_BUS <=  channel_threshold(3);
    when "011"    => ADC_THRESHOLD_BUS <=  channel_threshold(4);
    when "100"    => ADC_THRESHOLD_BUS <=  channel_threshold(5);
    when "101"    => ADC_THRESHOLD_BUS <=  channel_threshold(6);
    when "110"    => ADC_THRESHOLD_BUS <=  channel_threshold(7);
    when "111"    => ADC_THRESHOLD_BUS <=  channel_threshold(8);
  end case;
  end if;
--end if;
end process ADC_THRESHOLD_BUS_PROC;

ADC_IN_BUS_PROC: process (RESET, channel_counter)  begin
--if  rising_edge(CLOCK) then
  if (RESET = '1') then
  ADC_IN_BUS <= (others => '0');
  else
  case std_logic_vector(channel_counter(2 downto 0)) is
    when "000"    => ADC_IN_BUS <=  std_logic_vector(average(1))(9 downto 0);
    when "001"    => ADC_IN_BUS <=  std_logic_vector(average(2))(9 downto 0);
    when "010"    => ADC_IN_BUS <=  std_logic_vector(average(3))(9 downto 0);
    when "011"    => ADC_IN_BUS <=  std_logic_vector(average(4))(9 downto 0);
    when "100"    => ADC_IN_BUS <=  std_logic_vector(average(5))(9 downto 0);
    when "101"    => ADC_IN_BUS <=  std_logic_vector(average(6))(9 downto 0);
    when "110"    => ADC_IN_BUS <=  std_logic_vector(average(7))(9 downto 0);
    when "111"    => ADC_IN_BUS <=  std_logic_vector(average(8))(9 downto 0);
  end case;
  end if;
--end if;
end process ADC_IN_BUS_PROC;

SELECT_PEDESTAL_MEMORY_TO_READ: process(CLOCK) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    PED_DATA_OUT <= (others => '0');
  else    -- if TRB_PED_ADDR_IN(11 downto 8) = LOCAL_ID_IN then
    case TRB_PED_ADDR_IN(7 downto 5) is
      when "000" => PED_DATA_OUT <= channel_threshold(1)(15 downto 6);
      when "001" => PED_DATA_OUT <= channel_threshold(2)(15 downto 6);
      when "010" => PED_DATA_OUT <= channel_threshold(3)(15 downto 6);
      when "011" => PED_DATA_OUT <= channel_threshold(4)(15 downto 6);
      when "100" => PED_DATA_OUT <= channel_threshold(5)(15 downto 6);
      when "101" => PED_DATA_OUT <= channel_threshold(6)(15 downto 6);
      when "110" => PED_DATA_OUT <= channel_threshold(7)(15 downto 6);
      when "111" => PED_DATA_OUT <= channel_threshold(8)(15 downto 6);
    end case;
--  else
--    PED_DATA_OUT <= (others => 'Z');
  end if;
end if;
end process SELECT_PEDESTAL_MEMORY_TO_READ;

DELAYED_WRITE_ACK_PROCESS: process(RESET, CLOCK) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    delayed_write_ack <= (others => '0');
  else
    delayed_write_ack <= delayed_write_ack(1 downto 0) & PED_WRITE_IN;
  end if;
end if;
end process DELAYED_WRITE_ACK_PROCESS;
PED_WRITE_ACK_OUT        <= delayed_write_ack(2);

DELAYED_READ_ACK_PROCESS: process(RESET, CLOCK) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    delayed_read_ack <= (others => '0');
  else
    delayed_read_ack <= delayed_read_ack(1 downto 0) & PED_READ_IN;
  end if;
end if;
end process DELAYED_READ_ACK_PROCESS;
 PED_READ_ACK_OUT         <= delayed_read_ack(2); -- this line (read) is to be changed/removed after the output register is added to the RAM.

SELECT_PEDESTAL_MEMORY_TO_WRITE: process(RESET, CLOCK, PED_WRITE_IN, TRB_PED_ADDR_IN(2 downto 0), pedestal_calculation, acalcul_state) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    WRITE_PEDESTAL <= (others => '0');
  elsif PED_WRITE_IN = '1' then
      case TRB_PED_ADDR_IN(7 downto 5) is
        when "000" => WRITE_PEDESTAL <= "00000001";
        when "001" => WRITE_PEDESTAL <= "00000010";
        when "010" => WRITE_PEDESTAL <= "00000100";
        when "011" => WRITE_PEDESTAL <= "00001000";
        when "100" => WRITE_PEDESTAL <= "00010000";
        when "101" => WRITE_PEDESTAL <= "00100000";
        when "110" => WRITE_PEDESTAL <= "01000000";
        when "111" => WRITE_PEDESTAL <= "10000000";
      end case;
  elsif write_state = write_to_fifo then
      case std_logic_vector(channel_counter (2 downto 0) is
        when "000" => WRITE_PEDESTAL <= "00000001";
        when "001" => WRITE_PEDESTAL <= "00000010";
        when "010" => WRITE_PEDESTAL <= "00000100";
        when "011" => WRITE_PEDESTAL <= "00001000";
        when "100" => WRITE_PEDESTAL <= "00010000";
        when "101" => WRITE_PEDESTAL <= "00100000";
        when "110" => WRITE_PEDESTAL <= "01000000";
        when "111" => WRITE_PEDESTAL <= "10000000";
      end case;
  else
      WRITE_PEDESTAL <= (others => '0');
  end if;
end if;
end process SELECT_PEDESTAL_MEMORY_TO_WRITE;

NEXT_STATE_GEN: process(RESET, CLOCK) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    write_state <= idle;
    acalcul_state <= idle_ac;
  else
    write_state <= next_write_state;
    acalcul_state <= next_acalcul_state;
  end if;
end if;
end process NEXT_STATE_GEN;

DATA_VALID_PROCESS: process(RESET, CLOCK, write_state, pedestal_calculation) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    fee_data_write <= '0';
  else
      if (write_state = write_to_fifo) and pedestal_calculation = '0' then      --****************
        fee_data_write <= threshold_comparison_status(0);
      else
        fee_data_write <= '0';
      end if;
  end if;
end if;
end process DATA_VALID_PROCESS;

WRITE_RESULTS: process (RESET, write_state, sampling_end(5), channel_counter(3) )begin
  if(RESET = '1') then
    next_write_state <= idle;
  else
    case write_state is
    
      when IDLE       =>  if sampling_end(5) = '1' then
                      next_write_state <= wait_for_average;
                    else
                      next_write_state <= idle;
                    end if;
                
      when WAIT_FOR_AVERAGE =>  next_write_state <= wait_for_comparators;

      when WAIT_FOR_COMPARATORS => next_write_state <= wait_for_comp_status;

      when WAIT_FOR_COMP_STATUS => next_write_state <= write_to_fifo;

      when WRITE_TO_FIFO    =>  next_write_state <= test_completed; --inc_channel_counter;

--      when INC_CHANNEL_COUNTER  =>  next_write_state <= test_completed;
      
      when TEST_COMPLETED   =>  if channel_counter(3) = '1' then
                      next_write_state <= column_finished;
                    else
                      next_write_state <= write_to_fifo;
                    end if;

      when COLUMN_FINISHED  => next_write_state <= test_event_finished;

      when TEST_EVENT_FINISHED => if COLUMN_COUNTER(4 downto 0) = "00000" then
                      next_write_state <= event_finished_or_continue_pedestal;
                    else
                      next_write_state <= idle;
                    end if;
      when  event_finished_or_continue_pedestal => 
                    if pedestal_calculation = '1' then
                          if COLUMN_COUNTER(10 downto 5) = "000000" then
                                next_write_state <= send_out_thresholds;
                          else
                                next_write_state <= idle;
                          end if;
                    else
                        next_write_state <= event_finished;
                    end if;

      when EVENT_FINISHED   => next_write_state <= idle;

      when send_out_thresholds =>  next_write_state <= event_finished;

      when others       => next_write_state <= idle;

    end case;
  end if;
end process WRITE_RESULTS;

state_bits <=     x"0" when write_state = IDLE
               else x"1" when write_state = WAIT_FOR_AVERAGE
               else x"2" when write_state = WAIT_FOR_COMPARATORS
               else x"3" when write_state = WAIT_FOR_COMP_STATUS
               else x"4" when write_state = WRITE_TO_FIFO
               else x"5" when write_state = INC_CHANNEL_COUNTER
               else x"6" when write_state = TEST_COMPLETED
               else x"7" when write_state = COLUMN_FINISHED
               else x"8" when write_state = TEST_EVENT_FINISHED
               else x"9" when write_state = EVENT_FINISHED
               else x"F";
-- 
-- state_bits(0) <=  '0' when write_state = IDLE else '1';
-- state_bits(1) <= start_extended;
-- state_bits(2) <= ADC_RESULT_VALID;
-- state_bits(3) <= sampling_end(0);
-- 

SELECT_PEDESTAL_ADDRESS: process(RESET, CLOCK, write_state) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    PEDESTAL_ADDRESS <= (others => '0');
  else
    if write_state = idle then
      PEDESTAL_ADDRESS <= TRB_PED_ADDR_IN(4 downto 0);
    else 
      PEDESTAL_ADDRESS <= std_logic_vector(COLUMN_COUNTER(4 downto 0));
    end if;
  end if;
end if;
end process SELECT_PEDESTAL_ADDRESS;

ADVANCE_COLUMN_COUNTER: process(RESET, CLOCK, write_state) begin
if rising_edge(CLOCK) then
  if(RESET = '1') then
    COLUMN_COUNTER <= (others => '0');
  else
    if write_state = column_finished then
      COLUMN_COUNTER <= COLUMN_COUNTER + 1; -- "00001";
    end if;
  end if;
end if;
end process ADVANCE_COLUMN_COUNTER;

--********************** MK

  PEDESTAL_CALCULATION_PROC: process (RESET, acalcul_state, fee_trg_type, PEDESTAL_EVENT_COUNTER, sampling_end(7))begin
  if(RESET = '1') then
    next_acalcul_state <= idle_ac;
  else
    case acalcul_state is
    
      when idle_ac        =>  if pedestal_calculation = '1' and FEB_MUX_NEW_CHAN_RDY_IN = '1' then     --******************
                        next_acalcul_state <= first_pedestal_sample;
                      else
                        next_acalcul_state <= idle_ac;
                      end if;

      when first_pedestal_sample    =>  if sampling_end(7) = '1' then
                        next_acalcul_state <= write_ADC_to_memory;
                      else
                        next_acalcul_state <= first_pedestal_sample;
                      end if;

      when write_ADC_to_memory  => next_acalcul_state <= check_first_event_end;

      when check_first_event_end  => if COLUMN_COUNTER = "11111" then
                        next_acalcul_state <= wait_for_next_event;
                      else
                        next_acalcul_state <= synch_wait;
                      end if;
      when synch_wait       =>  if sampling_end(7) = '0' then
                        next_acalcul_state <= first_pedestal_sample;
                      else
                        next_acalcul_state <= synch_wait;
                      end if;

      when check_counter      =>  if PEDESTAL_EVENT_COUNTER = "111111" then
                        next_acalcul_state <= average_calcul_finished;
                      else
                        next_acalcul_state <= wait_for_next_event;
                      end if;

      when wait_for_next_event  => next_acalcul_state <= read_pedestal_value;   --*********????????????????????????

      when read_pedestal_value  => if sampling_end(7) = '1' then
                        next_acalcul_state <= sum_with_ADC;
                      else
                        next_acalcul_state <= read_pedestal_value;
                      end if;

      when sum_with_ADC     =>  next_acalcul_state <= write_sum_to_memory;

      when write_sum_to_memory  => next_acalcul_state <= check_ped_event_end;
      when check_ped_event_end  =>  if COLUMN_COUNTER = "11111" then
                        next_acalcul_state <= check_counter;
                      else
                        next_acalcul_state <= synch_wait_1;
                      end if;
      when synch_wait_1       =>  if sampling_end(7) = '0' then 
                        next_acalcul_state <= read_pedestal_value;
                      else
                        next_acalcul_state <= synch_wait_1;
                      end if;

      when average_calcul_finished => next_acalcul_state <= average_calcul_finished;
--      when average_calcul_finished => next_acalcul_state <= idle_ac;

      when others         => next_acalcul_state <= idle_ac;

    end case;
  end if;
end process PEDESTAL_CALCULATION_PROC;

end Behavioral;
